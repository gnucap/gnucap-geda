simulator language=verilog
// This File is part of gnucap-geda
// (C) 2012 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "asic" section

module PMOS_TRANSISTOR(D G S B);
// not yet
endmodule
hidemodule PMOS_TRANSISTOR

module NMOS_TRANSISTOR(D G S B);
// not yet
endmodule
hidemodule NMOS_TRANSISTOR

simulator lang=acs
