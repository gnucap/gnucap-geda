simulator language=verilog
// This File is part of gnucap-geda
// (C) 2012 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "switcap" section

module SWITCAP-capacitor(1 2);
// not yet.
endmodule
hidemodule SWITCAP-capacitor

simulator lang=acs
