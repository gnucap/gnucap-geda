simulator language=verilog
// This File is part of gnucap-geda
// (C) 2012 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "transistor" section

module BC547(1 2 3 4);
// nothing yet, just pins.
endmodule

simulator lang=acs
