simulator language=verilog
// This File is part of gnucap-geda
// (C) 2012 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "linear" section

// lm741-1.sym, missing pinseq=1,5?
module LM741(1 2 3 4 5 6 7);
// not yet
endmodule

module 555timer(1 2 3 4 5 6 7 8);
// not yet
endmodule

simulator lang=acs
