simulator language=verilog
// This File is part of gnucap-geda
// (C) 2015 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "74" section

module 7400(1 2 3);
// nothing yet
endmodule

module 7408(A B Y);
// nothing yet
endmodule

module 7432(A B Y);
// nothing yet
endmodule

module 7486(A B Y);
// nothing yet
endmodule

simulator lang=acs
