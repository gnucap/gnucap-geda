simulator language=verilog
// This File is part of gnucap-geda
// (C) 2012 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "connector" section

module HEADER3(1 2 3);
endmodule
hidemodule HEADER3

module DB25(SLCT,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25);
endmodule
hidemodule DB25

simulator lang=acs
