simulator language=verilog
// This File is part of gnucap-geda
// (C) 2015 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "74" section

module 7400(1 2 3);
// nothing yet
endmodule
hidemodule 7400

module 7408(A B Y);
// nothing yet
endmodule
hidemodule 7408

module 7432(A B Y);
// nothing yet
endmodule
hidemodule 7432

module 7486(A B Y);
// nothing yet
endmodule
hidemodule 7486

simulator lang=acs
