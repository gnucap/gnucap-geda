simulator language=verilog
// This File is part of gnucap-geda
// (C) 2015 Felix Salfelder
// GPLv3 or later

// mapping geda-symbols to actual devices
// "diode" section

module DIODE(1 2);
endmodule

module LEDseries(1 2);
endmodule

simulator lang=acs
